`include "tar_alu_sequence_item.sv"

`include "Alu_add_sequence.sv"
`include "Alu_sub_sequence.sv"
`include "Alu_and_sequence.sv"
`include "Alu_or_sequence.sv"
`include "Alu_xor_sequence.sv"
`include "Alu_undefined_opcode_sequence.sv"
`include "ALU_random_sequence.sv"
`include "tar_alu_sequencer.sv"
`include "tar_alu_driver.sv"
`include "tar_alu_monitor.sv"
`include "Alu_scoreboard.sv"
`include "subscriber.sv"
`include "alu_agent.sv"
`include "Alu_env.sv"